 

//------------------------------------------------------------------------------
// File       : and_gate.sv
// Author     : Punith R / 1BM24EC415
// Created    : 2026-02-08
// Module     : and_gate
// Project    : SystemVerilog and Verification (23EC6PE2SV)
// Faculty    : Prof. Ajaykumar Devarapalli
// Description: 2-input AND gate used for basic functional coverage example.
//------------------------------------------------------------------------------

module and_gate (
    input  logic a,
    input  logic b,
    output logic y
);

    assign y = a & b;

endmodule 
